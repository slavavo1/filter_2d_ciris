`define SIGNED_IN;
`define INTEL;
//`define FIFO_INTEL;